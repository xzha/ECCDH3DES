//$Id: mg78$
// Author: Nico Bellante
// nico@purdue.edu
// Lab Section: 337-03
// Description: Testbench for 3DES

`timescale 1ns / 1ps
module tb_des_TripleDES
(
);
	localparam NUM_BITS 		= 163; 	
	localparam NUM_INPUT_BITS 	= 3;
	localparam CLK_PERIOD 		= 3.33;
	localparam ROLLOVER_VAL 	= 10;
	localparam CHECK_DELAY 		= 1; // Check 1ns after the rising edge to allow for propagation delay

	parameter KEY_FILE 			= "./pythond3s/192bitkey.txt";
	parameter NUM_TEST_CASES    = 100;
	string IN_FILES [100] 		= {"./pythond3s/inputblock_0.txt", "./pythond3s/inputblock_1.txt", "./pythond3s/inputblock_2.txt", "./pythond3s/inputblock_3.txt", "./pythond3s/inputblock_4.txt", "./pythond3s/inputblock_5.txt", "./pythond3s/inputblock_6.txt", "./pythond3s/inputblock_7.txt", "./pythond3s/inputblock_8.txt", "./pythond3s/inputblock_9.txt", "./pythond3s/inputblock_10.txt", "./pythond3s/inputblock_11.txt", "./pythond3s/inputblock_12.txt", "./pythond3s/inputblock_13.txt", "./pythond3s/inputblock_14.txt", "./pythond3s/inputblock_15.txt", "./pythond3s/inputblock_16.txt", "./pythond3s/inputblock_17.txt", "./pythond3s/inputblock_18.txt", "./pythond3s/inputblock_19.txt", "./pythond3s/inputblock_20.txt", "./pythond3s/inputblock_21.txt", "./pythond3s/inputblock_22.txt", "./pythond3s/inputblock_23.txt", "./pythond3s/inputblock_24.txt", "./pythond3s/inputblock_25.txt", "./pythond3s/inputblock_26.txt", "./pythond3s/inputblock_27.txt", "./pythond3s/inputblock_28.txt", "./pythond3s/inputblock_29.txt", "./pythond3s/inputblock_30.txt", "./pythond3s/inputblock_31.txt", "./pythond3s/inputblock_32.txt", "./pythond3s/inputblock_33.txt", "./pythond3s/inputblock_34.txt", "./pythond3s/inputblock_35.txt", "./pythond3s/inputblock_36.txt", "./pythond3s/inputblock_37.txt", "./pythond3s/inputblock_38.txt", "./pythond3s/inputblock_39.txt", "./pythond3s/inputblock_40.txt", "./pythond3s/inputblock_41.txt", "./pythond3s/inputblock_42.txt", "./pythond3s/inputblock_43.txt", "./pythond3s/inputblock_44.txt", "./pythond3s/inputblock_45.txt", "./pythond3s/inputblock_46.txt", "./pythond3s/inputblock_47.txt", "./pythond3s/inputblock_48.txt", "./pythond3s/inputblock_49.txt", "./pythond3s/inputblock_50.txt", "./pythond3s/inputblock_51.txt", "./pythond3s/inputblock_52.txt", "./pythond3s/inputblock_53.txt", "./pythond3s/inputblock_54.txt", "./pythond3s/inputblock_55.txt", "./pythond3s/inputblock_56.txt", "./pythond3s/inputblock_57.txt", "./pythond3s/inputblock_58.txt", "./pythond3s/inputblock_59.txt", "./pythond3s/inputblock_60.txt", "./pythond3s/inputblock_61.txt", "./pythond3s/inputblock_62.txt", "./pythond3s/inputblock_63.txt", "./pythond3s/inputblock_64.txt", "./pythond3s/inputblock_65.txt", "./pythond3s/inputblock_66.txt", "./pythond3s/inputblock_67.txt", "./pythond3s/inputblock_68.txt", "./pythond3s/inputblock_69.txt", "./pythond3s/inputblock_70.txt", "./pythond3s/inputblock_71.txt", "./pythond3s/inputblock_72.txt", "./pythond3s/inputblock_73.txt", "./pythond3s/inputblock_74.txt", "./pythond3s/inputblock_75.txt", "./pythond3s/inputblock_76.txt", "./pythond3s/inputblock_77.txt", "./pythond3s/inputblock_78.txt", "./pythond3s/inputblock_79.txt", "./pythond3s/inputblock_80.txt", "./pythond3s/inputblock_81.txt", "./pythond3s/inputblock_82.txt", "./pythond3s/inputblock_83.txt", "./pythond3s/inputblock_84.txt", "./pythond3s/inputblock_85.txt", "./pythond3s/inputblock_86.txt", "./pythond3s/inputblock_87.txt", "./pythond3s/inputblock_88.txt", "./pythond3s/inputblock_89.txt", "./pythond3s/inputblock_90.txt", "./pythond3s/inputblock_91.txt", "./pythond3s/inputblock_92.txt", "./pythond3s/inputblock_93.txt", "./pythond3s/inputblock_94.txt", "./pythond3s/inputblock_95.txt", "./pythond3s/inputblock_96.txt", "./pythond3s/inputblock_97.txt", "./pythond3s/inputblock_98.txt", "./pythond3s/inputblock_99.txt"};	
	string OUT_FILES [100] 		= {"./pythond3s/outputofdes_0.txt", "./pythond3s/outputofdes_1.txt", "./pythond3s/outputofdes_2.txt", "./pythond3s/outputofdes_3.txt", "./pythond3s/outputofdes_4.txt", "./pythond3s/outputofdes_5.txt", "./pythond3s/outputofdes_6.txt", "./pythond3s/outputofdes_7.txt", "./pythond3s/outputofdes_8.txt", "./pythond3s/outputofdes_9.txt", "./pythond3s/outputofdes_10.txt", "./pythond3s/outputofdes_11.txt", "./pythond3s/outputofdes_12.txt", "./pythond3s/outputofdes_13.txt", "./pythond3s/outputofdes_14.txt", "./pythond3s/outputofdes_15.txt", "./pythond3s/outputofdes_16.txt", "./pythond3s/outputofdes_17.txt", "./pythond3s/outputofdes_18.txt", "./pythond3s/outputofdes_19.txt", "./pythond3s/outputofdes_20.txt", "./pythond3s/outputofdes_21.txt", "./pythond3s/outputofdes_22.txt", "./pythond3s/outputofdes_23.txt", "./pythond3s/outputofdes_24.txt", "./pythond3s/outputofdes_25.txt", "./pythond3s/outputofdes_26.txt", "./pythond3s/outputofdes_27.txt", "./pythond3s/outputofdes_28.txt", "./pythond3s/outputofdes_29.txt", "./pythond3s/outputofdes_30.txt", "./pythond3s/outputofdes_31.txt", "./pythond3s/outputofdes_32.txt", "./pythond3s/outputofdes_33.txt", "./pythond3s/outputofdes_34.txt", "./pythond3s/outputofdes_35.txt", "./pythond3s/outputofdes_36.txt", "./pythond3s/outputofdes_37.txt", "./pythond3s/outputofdes_38.txt", "./pythond3s/outputofdes_39.txt", "./pythond3s/outputofdes_40.txt", "./pythond3s/outputofdes_41.txt", "./pythond3s/outputofdes_42.txt", "./pythond3s/outputofdes_43.txt", "./pythond3s/outputofdes_44.txt", "./pythond3s/outputofdes_45.txt", "./pythond3s/outputofdes_46.txt", "./pythond3s/outputofdes_47.txt", "./pythond3s/outputofdes_48.txt", "./pythond3s/outputofdes_49.txt", "./pythond3s/outputofdes_50.txt", "./pythond3s/outputofdes_51.txt", "./pythond3s/outputofdes_52.txt", "./pythond3s/outputofdes_53.txt", "./pythond3s/outputofdes_54.txt", "./pythond3s/outputofdes_55.txt", "./pythond3s/outputofdes_56.txt", "./pythond3s/outputofdes_57.txt", "./pythond3s/outputofdes_58.txt", "./pythond3s/outputofdes_59.txt", "./pythond3s/outputofdes_60.txt", "./pythond3s/outputofdes_61.txt", "./pythond3s/outputofdes_62.txt", "./pythond3s/outputofdes_63.txt", "./pythond3s/outputofdes_64.txt", "./pythond3s/outputofdes_65.txt", "./pythond3s/outputofdes_66.txt", "./pythond3s/outputofdes_67.txt", "./pythond3s/outputofdes_68.txt", "./pythond3s/outputofdes_69.txt", "./pythond3s/outputofdes_70.txt", "./pythond3s/outputofdes_71.txt", "./pythond3s/outputofdes_72.txt", "./pythond3s/outputofdes_73.txt", "./pythond3s/outputofdes_74.txt", "./pythond3s/outputofdes_75.txt", "./pythond3s/outputofdes_76.txt", "./pythond3s/outputofdes_77.txt", "./pythond3s/outputofdes_78.txt", "./pythond3s/outputofdes_79.txt", "./pythond3s/outputofdes_80.txt", "./pythond3s/outputofdes_81.txt", "./pythond3s/outputofdes_82.txt", "./pythond3s/outputofdes_83.txt", "./pythond3s/outputofdes_84.txt", "./pythond3s/outputofdes_85.txt", "./pythond3s/outputofdes_86.txt", "./pythond3s/outputofdes_87.txt", "./pythond3s/outputofdes_88.txt", "./pythond3s/outputofdes_89.txt", "./pythond3s/outputofdes_90.txt", "./pythond3s/outputofdes_91.txt", "./pythond3s/outputofdes_92.txt", "./pythond3s/outputofdes_93.txt", "./pythond3s/outputofdes_94.txt", "./pythond3s/outputofdes_95.txt", "./pythond3s/outputofdes_96.txt", "./pythond3s/outputofdes_97.txt", "./pythond3s/outputofdes_98.txt", "./pythond3s/outputofdes_99.txt"};	
	integer i;
	integer j;
	integer key_f;
	integer out_f;
	integer in_block_f;

	integer current_test_case_index;
	integer verified_output_index = 0;

	// Declare test bench signals
	reg [0:63] tb_actual_input;
	reg [0:63] tb_actual_output;
	reg [0:NUM_TEST_CASES][0:7][7:0] tb_input_block;
	reg [0:NUM_TEST_CASES][0:7][7:0] tb_ciphertext_block;
	reg [0:23][7:0]tb_Sk;
	reg tb_data_valid_in;
	reg tb_data_valid_out;

	reg [0:NUM_TEST_CASES][0:7][7:0] tb_gold_ciphertext_3;

	reg tb_clk;
	reg tb_n_rst;


	// this task sends the input to the triple DES block with the proper data valid in and increments the index accordingly

	task input_data;
		input [0:63] data;
	begin
		@(negedge tb_clk);
		tb_data_valid_in = 1;
		tb_actual_input = data;
		@(posedge tb_clk);
		#(1);
		tb_data_valid_in = 0;
		current_test_case_index++;
	end
	endtask


	always
	begin
		tb_clk = 1'b0;
		#(CLK_PERIOD/2.0);
		tb_clk = 1'b1;
		#(CLK_PERIOD/2.0);
	end


	des_TripleDES DUTE(
		.input_block(tb_actual_input),
		.Sk          (tb_Sk),
		.is_encrypt  (1'b1),
		.clk         (tb_clk),
		.n_rst         (tb_n_rst),
		.data_valid_in (tb_data_valid_in),
		.data_valid_out(tb_data_valid_out),
		.output_block(tb_actual_output)
	);

	// this always block monitors the output of triple DES and checks if the output matches the correct output

	// !!! NOTE: if running in source, the posedge below must be changed to negedge !!! // 	

	always @ (posedge tb_clk)
	begin
		if (tb_data_valid_out == 1)
		begin
			assert(tb_actual_output == tb_gold_ciphertext_3[verified_output_index])
			begin
				$info("Everything looks good!");
			end
			else
			begin
				$error("UT OH! STUFF DOESNT LOOK RIGHT! ERRORROROROR!!!");
			end

			verified_output_index++;
		end
	end


	// Test bench process
	initial
	begin

		tb_data_valid_in = 1'b0;
		current_test_case_index = 0;
		
		/* this section will open the key file, input blocks, and correct output blocks 
		   the correct outputs will be used to verify it is encrypting properly */

		key_f = $fopen(KEY_FILE, "rb");

		for (i=0; i<24; i++)
		begin
			$fscanf(key_f,"%c",tb_Sk[i]);
		end
		
		$fclose(key_f);

		for (j=0; j<NUM_TEST_CASES; j++)
		begin

			in_block_f = $fopen(IN_FILES[j], "rb");
			out_f = $fopen(OUT_FILES[j], "rb");


			for (i=0; i<8; i++)
			begin
				$fscanf(out_f,"%c",tb_gold_ciphertext_3[j][i]);
				$fscanf(in_block_f,"%c",tb_input_block[j][i]);
			end

			$fclose(in_block_f);
			$fclose(out_f);

	    	end
		
		tb_n_rst = 1'b1;

		// Power-on Reset of the DUT
		#(0.1);
		tb_n_rst	= 1'b0; 	// Need to actually toggle this in order for it to actually run dependent always blocks
		#(CLK_PERIOD * 2.25);		// Release the reset away from a clock edge
		tb_n_rst	= 1'b1; 	// Deactivate the chip reset

		// Wait for a while to see normal operation
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);

		for (i=0; i<20; i++)
		begin
			input_data(tb_input_block[current_test_case_index]);
	    	end

		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
	
		input_data(tb_input_block[current_test_case_index]);
		input_data(tb_input_block[current_test_case_index]);

		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		
		input_data(tb_input_block[current_test_case_index]);
		
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);

		for (i=0; i<60; i++)
		begin
			input_data(tb_input_block[current_test_case_index]);
	    	end
		
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);
		#(CLK_PERIOD);

		input_data(tb_input_block[current_test_case_index]);


end

endmodule


// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);
// @(negedge tb_clk);

// 	assert(tb_gold_ciphertext_3 == tb_ciphertext_block)
// 	begin
// 		$info("Correct value!!!!!!!!!!!!!!!!!:D");
// 	end
// 	else
// 	begin
// 		$error("VALUES ARE NOT EQUAL!");
// 	end

// end




// 	// logic [63:0] tb_input_test_0 = 64'hee7da322ef81d7c5;
// 	// logic [63:0] tb_input_test_1 = 64'hefc4fb7e1ce98e4e;
// 	// logic [63:0] tb_input_test_2 = 64'he63ee286bfdc42fb;
// 	// logic [63:0] tb_input_test_3 = 64'hab4485038c80d0d3;
// 	// logic [63:0] tb_input_test_4 = 64'hc7d8cb57e75f832d;
// 	// logic [63:0] tb_input_test_5 = 64'hf84d0799d2035fed;
// 	// logic [63:0] tb_input_test_6 = 64'haccf25e223647a71;
// 	// logic [63:0] tb_input_test_7 = 64'hd3a27b14e23f52a6;
// 	// logic [63:0] tb_input_test_8 = 64'hfe23870431608e7d;
// 	// logic [63:0] tb_input_test_9 = 64'hbc620a9aa1efcce4;
// 	// logic [63:0] tb_input_test_10 = 64'hf0def6ffb307dbdc;
// 	// logic [63:0] tb_input_test_11 = 64'hba2eab4b42868c77;
// 	// logic [63:0] tb_input_test_12 = 64'ha7fd8505772ab14a;
// 	// logic [63:0] tb_input_test_13 = 64'ha880b2fe60349efb;
// 	// logic [63:0] tb_input_test_14 = 64'habc51d41aa40a92c;
// 	// logic [63:0] tb_input_test_15 = 64'hde63e9a4c56fb5db;
// 	// logic [63:0] tb_input_test_16 = 64'h812e8001d0a60e1e;
// 	// logic [63:0] tb_input_test_17 = 64'hd3e56e7980f3e649;
// 	// logic [63:0] tb_input_test_18 = 64'hc8a33802c862f4d1;
// 	// logic [63:0] tb_input_test_19 = 64'hee6496fb5b6916b8;
// 	// logic [63:0] tb_input_test_20 = 64'h81fecd943d72a8b3;
// 	// logic [63:0] tb_input_test_21 = 64'hd5b1a23ff6d7c73b;
// 	// logic [63:0] tb_input_test_22 = 64'hff1005ecd13e41b4;
// 	// logic [63:0] tb_input_test_23 = 64'hcc99a205c65e4f69;
// 	// logic [63:0] tb_input_test_24 = 64'hf792b2b128984be4;
// 	// logic [63:0] tb_input_test_25 = 64'had59fc90391eb101;
// 	// logic [63:0] tb_input_test_26 = 64'hc5e6b52ac4bffc55;
// 	// logic [63:0] tb_input_test_27 = 64'hc68a9fb45da7462d;
// 	// logic [63:0] tb_input_test_28 = 64'h80e54c355722d5e9;
// 	// logic [63:0] tb_input_test_29 = 64'he587b24599ce3b2f;
// 	// logic [63:0] tb_input_test_30 = 64'hd6604e34aadd00b4;
// 	// logic [63:0] tb_input_test_31 = 64'hbe9b95aa4005cac7;
// 	// logic [63:0] tb_input_test_32 = 64'hf62c032e9d176052;
// 	// logic [63:0] tb_input_test_33 = 64'ha377758f6508eac3;
// 	// logic [63:0] tb_input_test_34 = 64'hde32cb4fc3145ba6;
// 	// logic [63:0] tb_input_test_35 = 64'hb3e10e816cacb555;
// 	// logic [63:0] tb_input_test_36 = 64'h83935e8d99c8acfe;
// 	// logic [63:0] tb_input_test_37 = 64'hd088c203239e4d3c;
// 	// logic [63:0] tb_input_test_38 = 64'hd127b03978fde75c;
// 	// logic [63:0] tb_input_test_39 = 64'h96de06c1049c3e27;
// 	// logic [63:0] tb_input_test_40 = 64'ha352a03dc1f019d4;
// 	// logic [63:0] tb_input_test_41 = 64'hf815dfafad802886;
// 	// logic [63:0] tb_input_test_42 = 64'h84fa63122be1832f;
// 	// logic [63:0] tb_input_test_43 = 64'hfc92c004b7345c2a;
// 	// logic [63:0] tb_input_test_44 = 64'hc57e0ac95be682ee;
// 	// logic [63:0] tb_input_test_45 = 64'ha88bdb6d22d0f550;
// 	// logic [63:0] tb_input_test_46 = 64'haf2e9fea6f8ca50b;
// 	// logic [63:0] tb_input_test_47 = 64'ha792403806d276cc;
// 	// logic [63:0] tb_input_test_48 = 64'haef63c68797702a6;
// 	// logic [63:0] tb_input_test_49 = 64'h896ef4c1ad7c337b;
// 	// logic [63:0] tb_input_test_50 = 64'hdc46080119023b7e;
// 	// logic [63:0] tb_input_test_51 = 64'hae374c7c474a6080;
// 	// logic [63:0] tb_input_test_52 = 64'hbe2d76d3e726ffbb;
// 	// logic [63:0] tb_input_test_53 = 64'hc6211d71f533abda;
// 	// logic [63:0] tb_input_test_54 = 64'ha750aeeec9f3a5e5;
// 	// logic [63:0] tb_input_test_55 = 64'hb6241026d286280e;
// 	// logic [63:0] tb_input_test_56 = 64'hb76d5de0dddd3ea4;
// 	// logic [63:0] tb_input_test_57 = 64'h9fafda0b24d47bd1;
// 	// logic [63:0] tb_input_test_58 = 64'he28852bc6c5b280c;
// 	// logic [63:0] tb_input_test_59 = 64'hf43e408d8a100651;
// 	// logic [63:0] tb_input_test_60 = 64'h84e5583e3dd5cf4d;
// 	// logic [63:0] tb_input_test_61 = 64'h9c112b6097c2f355;
// 	// logic [63:0] tb_input_test_62 = 64'hc60fbcd38168fc74;
// 	// logic [63:0] tb_input_test_63 = 64'h8bee811784185829;
// 	// logic [63:0] tb_input_test_64 = 64'hc8d86dee9ccd15b0;
// 	// logic [63:0] tb_input_test_65 = 64'h98be7e8e754089e5;
// 	// logic [63:0] tb_input_test_66 = 64'hbb54298a80c804bc;
// 	// logic [63:0] tb_input_test_67 = 64'he613729868035c0e;
// 	// logic [63:0] tb_input_test_68 = 64'h8ad16a04e26e096f;
// 	// logic [63:0] tb_input_test_69 = 64'hbbc1ae75e97f6ca2;
// 	// logic [63:0] tb_input_test_70 = 64'hfd6fb8d151103f43;
// 	// logic [63:0] tb_input_test_71 = 64'hf09cc2631a5e1a28;
// 	// logic [63:0] tb_input_test_72 = 64'he3d85fed95860f77;
// 	// logic [63:0] tb_input_test_73 = 64'hc8d1ff10b9127ac6;
// 	// logic [63:0] tb_input_test_74 = 64'hcfd032dd60275355;
// 	// logic [63:0] tb_input_test_75 = 64'hf95ed35f2c149e57;
// 	// logic [63:0] tb_input_test_76 = 64'hae43825527b49ac6;
// 	// logic [63:0] tb_input_test_77 = 64'haae9d158af0ab0e0;
// 	// logic [63:0] tb_input_test_78 = 64'hb8057817ec9897ec;
// 	// logic [63:0] tb_input_test_79 = 64'hdcfa4200c688675b;
// 	// logic [63:0] tb_input_test_80 = 64'hb97ff3281d464035;
// 	// logic [63:0] tb_input_test_81 = 64'he05883bfbf868702;
// 	// logic [63:0] tb_input_test_82 = 64'hb9140ab0f6ea935e;
// 	// logic [63:0] tb_input_test_83 = 64'he149fd9cdc507cf0;
// 	// logic [63:0] tb_input_test_84 = 64'h91bff05713446337;
// 	// logic [63:0] tb_input_test_85 = 64'he34dd73ed588f8a8;
// 	// logic [63:0] tb_input_test_86 = 64'haaeba9b6beaf761e;
// 	// logic [63:0] tb_input_test_87 = 64'hd44a5bef1fc25a44;
// 	// logic [63:0] tb_input_test_88 = 64'hb0b8d039d2124881;
// 	// logic [63:0] tb_input_test_89 = 64'h867cef9aa48188e9;
// 	// logic [63:0] tb_input_test_90 = 64'haaf52b18a4d75398;
// 	// logic [63:0] tb_input_test_91 = 64'hc7d0749f7ca9bdc9;
// 	// logic [63:0] tb_input_test_92 = 64'hae105c72b4928192;
// 	// logic [63:0] tb_input_test_93 = 64'he04c679c633dbf88;
// 	// logic [63:0] tb_input_test_94 = 64'he3a0d6c0c020fe26;
// 	// logic [63:0] tb_input_test_95 = 64'hbccb52a761358cd2;
// 	// logic [63:0] tb_input_test_96 = 64'ha00d585e88e7c347;
// 	// logic [63:0] tb_input_test_97 = 64'hca9ffe8a52ce99fa;
// 	// logic [63:0] tb_input_test_98 = 64'he0654887d862b2ab;
// 	// logic [63:0] tb_input_test_99 = 64'h9904f4dddfcddb83;
// 	// logic [63:0] tb_input_test_100 = 64'hefe1f5fbcb0042ac;
// 	// logic [63:0] tb_input_test_101 = 64'hb41a84b490afa9f4;
// 	// logic [63:0] tb_input_test_102 = 64'ha1dad8dc3e981deb;
// 	// logic [63:0] tb_input_test_103 = 64'h9424d52e16c8cbcb;
// 	// logic [63:0] tb_input_test_104 = 64'haaa279bb2a44e756;
// 	// logic [63:0] tb_input_test_105 = 64'he228b73f39450da9;
// 	// logic [63:0] tb_input_test_106 = 64'he76eb611c5f8c11f;
// 	// logic [63:0] tb_input_test_107 = 64'hc96ab2077c918084;
// 	// logic [63:0] tb_input_test_108 = 64'hef190972271d71d7;
// 	// logic [63:0] tb_input_test_109 = 64'ha7f0907fc0c98e72;
// 	// logic [63:0] tb_input_test_110 = 64'hc12352a99593c974;
// 	// logic [63:0] tb_input_test_111 = 64'h9c2138ace1715734;
// 	// logic [63:0] tb_input_test_112 = 64'h9e112964176bef06;
// 	// logic [63:0] tb_input_test_113 = 64'hf141f70ce5f17618;
// 	// logic [63:0] tb_input_test_114 = 64'ha96f58c74a0f8097;
// 	// logic [63:0] tb_input_test_115 = 64'hffd6a24dc727dc3b;
// 	// logic [63:0] tb_input_test_116 = 64'h92fc0960f0313fc6;
// 	// logic [63:0] tb_input_test_117 = 64'hed3881eece9627fc;
// 	// logic [63:0] tb_input_test_118 = 64'he6d48b6b873738ab;
// 	// logic [63:0] tb_input_test_119 = 64'h9df74f4c543e54c4;
// 	// logic [63:0] tb_input_test_120 = 64'he482c862c2c5ce02;
// 	// logic [63:0] tb_input_test_121 = 64'hb30e8f7d6d1619a3;
// 	// logic [63:0] tb_input_test_122 = 64'h9ff1d99b6a38c654;
// 	// logic [63:0] tb_input_test_123 = 64'hb5e40bf78495f8cb;
// 	// logic [63:0] tb_input_test_124 = 64'hdda70efe9c4f5907;
// 	// logic [63:0] tb_input_test_125 = 64'hf311cf1cd4379666;
// 	// logic [63:0] tb_input_test_126 = 64'hcba66d434b473ab9;
// 	// logic [63:0] tb_input_test_127 = 64'h8b9e29cc6626c303;
// 	// logic [63:0] tb_input_test_128 = 64'hbafc5f44aa415831;
// 	// logic [63:0] tb_input_test_129 = 64'h9a3244bd8ed91243;
// 	// logic [63:0] tb_input_test_130 = 64'hada631206af6f394;
// 	// logic [63:0] tb_input_test_131 = 64'hd6082f24ab802c34;
// 	// logic [63:0] tb_input_test_132 = 64'h813cd61e0bd1adee;
// 	// logic [63:0] tb_input_test_133 = 64'hcaf02d015da3e2f4;
// 	// logic [63:0] tb_input_test_134 = 64'h99eabf8865f7dcf9;
// 	// logic [63:0] tb_input_test_135 = 64'h8edba82b50cfe841;
// 	// logic [63:0] tb_input_test_136 = 64'heff3a7dfb9acd522;
// 	// logic [63:0] tb_input_test_137 = 64'h8fac6ad6949d73e8;
// 	// logic [63:0] tb_input_test_138 = 64'h91c1fad98942b1b8;
// 	// logic [63:0] tb_input_test_139 = 64'h8fb6141b1a614801;
// 	// logic [63:0] tb_input_test_140 = 64'hedd622e01d3e139e;
// 	// logic [63:0] tb_input_test_141 = 64'he2600aae943e2e92;
// 	// logic [63:0] tb_input_test_142 = 64'ha39a452e543c9d16;
// 	// logic [63:0] tb_input_test_143 = 64'hd58c52bac9398bba;
// 	// logic [63:0] tb_input_test_144 = 64'hcf867c2a1814a095;
// 	// logic [63:0] tb_input_test_145 = 64'hf9b466a9be74f436;
// 	// logic [63:0] tb_input_test_146 = 64'he60951879ece2f3b;
// 	// logic [63:0] tb_input_test_147 = 64'hf8d3e21c0422f0e1;
// 	// logic [63:0] tb_input_test_148 = 64'he1e703bf586f7780;
// 	// logic [63:0] tb_input_test_149 = 64'hd347bf6ad86722a5;
// 	// logic [63:0] tb_input_test_150 = 64'hc7ee5523505a4922;
// 	// logic [63:0] tb_input_test_151 = 64'hcb2d53e29f17acd6;
// 	// logic [63:0] tb_input_test_152 = 64'hfe7d710646e542b6;
// 	// logic [63:0] tb_input_test_153 = 64'hca18683c18720758;
// 	// logic [63:0] tb_input_test_154 = 64'hf4c56db0988985f4;
// 	// logic [63:0] tb_input_test_155 = 64'hf1738f27528bb870;
// 	// logic [63:0] tb_input_test_156 = 64'he48e486aa511efa6;
// 	// logic [63:0] tb_input_test_157 = 64'hd997e315681beded;
// 	// logic [63:0] tb_input_test_158 = 64'hbdda2661eb242495;
// 	// logic [63:0] tb_input_test_159 = 64'he8fd70c9974d0170;
// 	// logic [63:0] tb_input_test_160 = 64'hd4695cf26a9608bb;
// 	// logic [63:0] tb_input_test_161 = 64'hda377d88346e0b38;
// 	// logic [63:0] tb_input_test_162 = 64'hc49e4b4d3b1786ad;
// 	// logic [63:0] tb_input_test_163 = 64'hd2be5d9c46669d72;
// 	// logic [63:0] tb_input_test_164 = 64'hda1db9fc06e05c6c;
// 	// logic [63:0] tb_input_test_165 = 64'hd2de40832ea08c1a;
// 	// logic [63:0] tb_input_test_166 = 64'hcef83175210c09d2;
// 	// logic [63:0] tb_input_test_167 = 64'hf6f6f20605729020;
// 	// logic [63:0] tb_input_test_168 = 64'hce17ea57e161c1a4;
// 	// logic [63:0] tb_input_test_169 = 64'h82b8e7eb940f4720;
// 	// logic [63:0] tb_input_test_170 = 64'hdb32c09ec3ac7a3b;
// 	// logic [63:0] tb_input_test_171 = 64'hbb7003fb972a7f6d;
// 	// logic [63:0] tb_input_test_172 = 64'hcb78289a0ab146c0;
// 	// logic [63:0] tb_input_test_173 = 64'hb1340588cd7debff;
// 	// logic [63:0] tb_input_test_174 = 64'hdf39876324d3457a;
// 	// logic [63:0] tb_input_test_175 = 64'hdae691cc003118b1;
// 	// logic [63:0] tb_input_test_176 = 64'hda64f92d68f034e4;
// 	// logic [63:0] tb_input_test_177 = 64'hc56b72f060d3cf2e;
// 	// logic [63:0] tb_input_test_178 = 64'hb251842d9aa6016c;
// 	// logic [63:0] tb_input_test_179 = 64'hd162edf4a2fb0a48;
// 	// logic [63:0] tb_input_test_180 = 64'headc1fba95ace08d;
// 	// logic [63:0] tb_input_test_181 = 64'ha8b0c00150950be4;
// 	// logic [63:0] tb_input_test_182 = 64'hfcd33f8fae6125c5;
// 	// logic [63:0] tb_input_test_183 = 64'h9cec4b93217104c1;
// 	// logic [63:0] tb_input_test_184 = 64'hc2b0e5811c3e9322;
// 	// logic [63:0] tb_input_test_185 = 64'h96466e14b40edb51;
// 	// logic [63:0] tb_input_test_186 = 64'h9da67f24d6d589ea;
// 	// logic [63:0] tb_input_test_187 = 64'h89819312f2832cd9;
// 	// logic [63:0] tb_input_test_188 = 64'hbf7acba64f69cba7;
// 	// logic [63:0] tb_input_test_189 = 64'h82104a03c57ed2b9;
// 	// logic [63:0] tb_input_test_190 = 64'hd288bf2ef6dd5a0d;
// 	// logic [63:0] tb_input_test_191 = 64'ha71c6d70bed8efd0;
// 	// logic [63:0] tb_input_test_192 = 64'h9b2787323f53f0d1;
// 	// logic [63:0] tb_input_test_193 = 64'hc7d17603de97795f;
// 	// logic [63:0] tb_input_test_194 = 64'hf403d88c32b5a35d;
// 	// logic [63:0] tb_input_test_195 = 64'hf9985f2b43d95f54;
// 	// logic [63:0] tb_input_test_196 = 64'hfeb53640c2f2823b;
// 	// logic [63:0] tb_input_test_197 = 64'h9d5580fdbdd67839;
// 	// logic [63:0] tb_input_test_198 = 64'hfe516bb05343f590;
// 	// logic [63:0] tb_input_test_199 = 64'had7b4812fe2b75b4;
// 	// logic [63:0] tb_input_test_200 = 64'h8196810b1fc10c9d;
// 	// logic [63:0] tb_input_test_201 = 64'hb71e2b8aedef89eb;
// 	// logic [63:0] tb_input_test_202 = 64'h998d0e9949f522e0;
// 	// logic [63:0] tb_input_test_203 = 64'h93dde0aff7452886;
// 	// logic [63:0] tb_input_test_204 = 64'hea3b4e10ff08aab0;
// 	// logic [63:0] tb_input_test_205 = 64'h89069632c8cb6c4f;
// 	// logic [63:0] tb_input_test_206 = 64'h855ef3f69189625d;
// 	// logic [63:0] tb_input_test_207 = 64'h84f4b6a9a60973f1;
// 	// logic [63:0] tb_input_test_208 = 64'h8ceb634bb48499ab;
// 	// logic [63:0] tb_input_test_209 = 64'hc76a712c85f4e65a;
// 	// logic [63:0] tb_input_test_210 = 64'hfd3a397b5c87cbab;
// 	// logic [63:0] tb_input_test_211 = 64'h944cce5690073cbc;
// 	// logic [63:0] tb_input_test_212 = 64'h98808c0a0d6e5368;
// 	// logic [63:0] tb_input_test_213 = 64'he90233cbf2460c8d;
// 	// logic [63:0] tb_input_test_214 = 64'ha1a0768bd0f53228;
// 	// logic [63:0] tb_input_test_215 = 64'hd0fbfba26ae2d5c5;
// 	// logic [63:0] tb_input_test_216 = 64'ha1ef0a4be85fa4be;
// 	// logic [63:0] tb_input_test_217 = 64'h8105fda61644c856;
// 	// logic [63:0] tb_input_test_218 = 64'h881082a053551b7c;
// 	// logic [63:0] tb_input_test_219 = 64'h8e3fd007259ba28b;
// 	// logic [63:0] tb_input_test_220 = 64'hdad728328af1d600;
// 	// logic [63:0] tb_input_test_221 = 64'h92f764b97031a585;
// 	// logic [63:0] tb_input_test_222 = 64'he78818111839fa48;
// 	// logic [63:0] tb_input_test_223 = 64'h9a830d42e8b2df3e;
// 	// logic [63:0] tb_input_test_224 = 64'hf14a88b7c58874d7;
// 	// logic [63:0] tb_input_test_225 = 64'hf2892af4b40bdc68;
// 	// logic [63:0] tb_input_test_226 = 64'h8b4fc7266b504997;
// 	// logic [63:0] tb_input_test_227 = 64'h90f9e1c196531c57;
// 	// logic [63:0] tb_input_test_228 = 64'hc5a06586e45ff9c1;
// 	// logic [63:0] tb_input_test_229 = 64'ha0944ab2a205c9c3;
// 	// logic [63:0] tb_input_test_230 = 64'hfab578f2759e52ab;
// 	// logic [63:0] tb_input_test_231 = 64'h9357b9aad06b0218;
// 	// logic [63:0] tb_input_test_232 = 64'h860f1712efe91f94;
// 	// logic [63:0] tb_input_test_233 = 64'hba89d8d2aa102352;
// 	// logic [63:0] tb_input_test_234 = 64'hc55c1c606c293c99;
// 	// logic [63:0] tb_input_test_235 = 64'he9f76ffbc7181f60;
// 	// logic [63:0] tb_input_test_236 = 64'hd844813d7f21bc41;
// 	// logic [63:0] tb_input_test_237 = 64'hb2093552eb4f49ed;
// 	// logic [63:0] tb_input_test_238 = 64'hdf0e8c643f60f386;
// 	// logic [63:0] tb_input_test_239 = 64'hf20048bf02dc4c22;
// 	// logic [63:0] tb_input_test_240 = 64'h9b3e1a0a8016ecf6;
// 	// logic [63:0] tb_input_test_241 = 64'he4b7e5476b6c94f4;
// 	// logic [63:0] tb_input_test_242 = 64'hcfcacdc1aa0c6c29;
// 	// logic [63:0] tb_input_test_243 = 64'hf255bf406e9ca984;
// 	// logic [63:0] tb_input_test_244 = 64'ha6923205be5f235d;
// 	// logic [63:0] tb_input_test_245 = 64'hcc502d86f2d2333b;
// 	// logic [63:0] tb_input_test_246 = 64'hd6b76d36ace2a3d7;
// 	// logic [63:0] tb_input_test_247 = 64'h9e7923c57b3c54ea;
// 	// logic [63:0] tb_input_test_248 = 64'h90491249158e29aa;
// 	// logic [63:0] tb_input_test_249 = 64'haa7531300753dbc1;
// 	// logic [63:0] tb_input_test_250 = 64'h98cc4c83d770d05e;
// 	// logic [63:0] tb_input_test_251 = 64'hce789a643d2bbfc5;
// 	// logic [63:0] tb_input_test_252 = 64'hf7926f082479a98b;
// 	// logic [63:0] tb_input_test_253 = 64'haf57fd4458a26467;
// 	// logic [63:0] tb_input_test_254 = 64'ha95da027b2ad8042;
// 	// logic [63:0] tb_input_test_255 = 64'hbd21f799c6f54ee3;
// 	// logic [63:0] tb_input_test_256 = 64'hf05a2eb4792f083f;
// 	// logic [63:0] tb_input_test_257 = 64'hd7a083335b3b273e;
// 	// logic [63:0] tb_input_test_258 = 64'hebba85cda4cb00e7;
// 	// logic [63:0] tb_input_test_259 = 64'hd34f81807dec03f7;
// 	// logic [63:0] tb_input_test_260 = 64'hdf6c8410f44e8686;
// 	// logic [63:0] tb_input_test_261 = 64'hd3563c46e2cae1f3;
// 	// logic [63:0] tb_input_test_262 = 64'hb92ac7e730499a36;
// 	// logic [63:0] tb_input_test_263 = 64'hefc9cf8c3496b742;
// 	// logic [63:0] tb_input_test_264 = 64'hd1fddb3670481b20;
// 	// logic [63:0] tb_input_test_265 = 64'h95d4388c91821b49;
// 	// logic [63:0] tb_input_test_266 = 64'h9570c05de62b985f;
// 	// logic [63:0] tb_input_test_267 = 64'hc9b1065cd66b4cb1;
// 	// logic [63:0] tb_input_test_268 = 64'ha9a6c758a7aabb53;
// 	// logic [63:0] tb_input_test_269 = 64'hff25d0ce9a012fc5;
// 	// logic [63:0] tb_input_test_270 = 64'hf86c56942fcc9880;
// 	// logic [63:0] tb_input_test_271 = 64'hecb8f5a2607b113d;
// 	// logic [63:0] tb_input_test_272 = 64'haaa33cd855054a60;
// 	// logic [63:0] tb_input_test_273 = 64'hc42af4bcf0fc1077;
// 	// logic [63:0] tb_input_test_274 = 64'hf8a6ff456474edd7;
// 	// logic [63:0] tb_input_test_275 = 64'h8234e6e3ab495632;
// 	// logic [63:0] tb_input_test_276 = 64'h886ad407208e76dc;
// 	// logic [63:0] tb_input_test_277 = 64'h97efd22aecbba7c8;
// 	// logic [63:0] tb_input_test_278 = 64'hc218253b5d11a973;
// 	// logic [63:0] tb_input_test_279 = 64'hebb0d847843d9752;
// 	// logic [63:0] tb_input_test_280 = 64'hc0b8d1e457fb5aad;
// 	// logic [63:0] tb_input_test_281 = 64'h8313c3b33924e603;
// 	// logic [63:0] tb_input_test_282 = 64'h9b00e231bca94657;
// 	// logic [63:0] tb_input_test_283 = 64'hfd81cf45b924e469;
// 	// logic [63:0] tb_input_test_284 = 64'hc389bd9247c38f17;
// 	// logic [63:0] tb_input_test_285 = 64'h8584054488c20158;
// 	// logic [63:0] tb_input_test_286 = 64'hf727995677ff9f98;
// 	// logic [63:0] tb_input_test_287 = 64'hdaf08a822bdf851d;
// 	// logic [63:0] tb_input_test_288 = 64'hea1aa727188a8669;
// 	// logic [63:0] tb_input_test_289 = 64'hf052a4074208de24;
// 	// logic [63:0] tb_input_test_290 = 64'hd51cc98c785d6385;
// 	// logic [63:0] tb_input_test_291 = 64'hc7a1307876437572;
// 	// logic [63:0] tb_input_test_292 = 64'hb6bf7b8e13af1f4e;
// 	// logic [63:0] tb_input_test_293 = 64'he79ff5a0d7683e43;
// 	// logic [63:0] tb_input_test_294 = 64'hc130bf272fe5e128;
// 	// logic [63:0] tb_input_test_295 = 64'ha699ff0ec428e44a;
// 	// logic [63:0] tb_input_test_296 = 64'ha7b62cdda938c1df;
// 	// logic [63:0] tb_input_test_297 = 64'h882d45f79f3cf782;
// 	// logic [63:0] tb_input_test_298 = 64'hffad8812b13f623f;
// 	// logic [63:0] tb_input_test_299 = 64'hd4d48c645af5e4e7;
// 	// logic [63:0] tb_input_test_300 = 64'hf470953dce93047a;
// 	// logic [63:0] tb_input_test_301 = 64'hb07180f98bf80882;
// 	// logic [63:0] tb_input_test_302 = 64'hc9779f22d4732050;
// 	// logic [63:0] tb_input_test_303 = 64'hb2c05840d934a76b;
// 	// logic [63:0] tb_input_test_304 = 64'hb7d12f85a3b5b831;
// 	// logic [63:0] tb_input_test_305 = 64'hd0013cd9601183f2;
// 	// logic [63:0] tb_input_test_306 = 64'h81591524e577e957;
// 	// logic [63:0] tb_input_test_307 = 64'haf29a190f7d8a259;
// 	// logic [63:0] tb_input_test_308 = 64'hd628d2370912981b;
// 	// logic [63:0] tb_input_test_309 = 64'hab9e81a3157b05fc;
// 	// logic [63:0] tb_input_test_310 = 64'haa186a428d5bb096;
// 	// logic [63:0] tb_input_test_311 = 64'hcbcde2126572dcda;
// 	// logic [63:0] tb_input_test_312 = 64'hba803e38a206c63e;
// 	// logic [63:0] tb_input_test_313 = 64'hd20894bb394f1013;
// 	// logic [63:0] tb_input_test_314 = 64'hb9e796ae366af9ed;
// 	// logic [63:0] tb_input_test_315 = 64'hc42631cc7e228657;
// 	// logic [63:0] tb_input_test_316 = 64'ha833a3be28304d85;
// 	// logic [63:0] tb_input_test_317 = 64'hadd54af0c38d6525;
// 	// logic [63:0] tb_input_test_318 = 64'hd1ebc6d6edfc4e67;
// 	// logic [63:0] tb_input_test_319 = 64'ha1b2918b23a915ab;
// 	// logic [63:0] tb_input_test_320 = 64'h9fd5b6adc0fbb3a4;
// 	// logic [63:0] tb_input_test_321 = 64'hea9dfab9ad64c43a;
// 	// logic [63:0] tb_input_test_322 = 64'hd0dce82105a0868b;
// 	// logic [63:0] tb_input_test_323 = 64'hf86a04f91838a7e3;
// 	// logic [63:0] tb_input_test_324 = 64'h98406e2225cfc050;
// 	// logic [63:0] tb_input_test_325 = 64'hd7a9d8e95397803e;
// 	// logic [63:0] tb_input_test_326 = 64'he3dbbbe339303f3e;
// 	// logic [63:0] tb_input_test_327 = 64'h97171666b52dc735;
// 	// logic [63:0] tb_input_test_328 = 64'h8764c6fd476d6b93;
// 	// logic [63:0] tb_input_test_329 = 64'hbef741536ca26d5d;
// 	// logic [63:0] tb_input_test_330 = 64'h99dcaf7371cc3d29;
// 	// logic [63:0] tb_input_test_331 = 64'hee984f20e3f300c5;
// 	// logic [63:0] tb_input_test_332 = 64'hd835fd2127618560;
// 	// logic [63:0] tb_input_test_333 = 64'h8b863fd8f1f5faba;
// 	// logic [63:0] tb_input_test_334 = 64'hef42ff7ed5319741;
// 	// logic [63:0] tb_input_test_335 = 64'h995b4bf7df798c9b;
// 	// logic [63:0] tb_input_test_336 = 64'h9f4abd60b3c6ddb7;
// 	// logic [63:0] tb_input_test_337 = 64'h9a736d0ce7de57d3;
// 	// logic [63:0] tb_input_test_338 = 64'ha0d19515d513af5b;
// 	// logic [63:0] tb_input_test_339 = 64'hc81b1a18b422f96a;
// 	// logic [63:0] tb_input_test_340 = 64'hbbcc537da8720cb7;
// 	// logic [63:0] tb_input_test_341 = 64'ha02678826286bd3f;
// 	// logic [63:0] tb_input_test_342 = 64'h9c6039152f52514b;
// 	// logic [63:0] tb_input_test_343 = 64'h8926ba6891751383;
// 	// logic [63:0] tb_input_test_344 = 64'he6d016192da53be5;
// 	// logic [63:0] tb_input_test_345 = 64'h849de190642426f8;
// 	// logic [63:0] tb_input_test_346 = 64'h8fca6a78fa335b0c;
// 	// logic [63:0] tb_input_test_347 = 64'hdf26eeda27e10709;
// 	// logic [63:0] tb_input_test_348 = 64'haadea17c1cb2bdbc;
// 	// logic [63:0] tb_input_test_349 = 64'hb79dd0ff61abbcec;
// 	// logic [63:0] tb_input_test_350 = 64'h9a9bbda60a61ff8e;
// 	// logic [63:0] tb_input_test_351 = 64'hd4f0478a5ca392d1;
// 	// logic [63:0] tb_input_test_352 = 64'h9458eafde4268a42;
// 	// logic [63:0] tb_input_test_353 = 64'h9e25ce4edeb5a0a3;
// 	// logic [63:0] tb_input_test_354 = 64'ha3c8fa4caafe8691;
// 	// logic [63:0] tb_input_test_355 = 64'hd18787a8965ea317;
// 	// logic [63:0] tb_input_test_356 = 64'h917e45eb91ffa21c;
// 	// logic [63:0] tb_input_test_357 = 64'hff6ee7d2fb5c2556;
// 	// logic [63:0] tb_input_test_358 = 64'hdc02317617909bec;
// 	// logic [63:0] tb_input_test_359 = 64'h8b5a553d993d4f28;
// 	// logic [63:0] tb_input_test_360 = 64'ha0c69c34c71f5749;
// 	// logic [63:0] tb_input_test_361 = 64'h8020d041c76c8b76;
// 	// logic [63:0] tb_input_test_362 = 64'ha3917abaf4aa1e66;
// 	// logic [63:0] tb_input_test_363 = 64'hfb43af8a17b817d8;
// 	// logic [63:0] tb_input_test_364 = 64'h9f7bd89b23324049;
// 	// logic [63:0] tb_input_test_365 = 64'hf27d208aaf3e509b;
// 	// logic [63:0] tb_input_test_366 = 64'h9da9ee16f7866a6e;
// 	// logic [63:0] tb_input_test_367 = 64'hd2d7162794840329;
// 	// logic [63:0] tb_input_test_368 = 64'hb13aea857229b43a;
// 	// logic [63:0] tb_input_test_369 = 64'hbd52f0a6d625f619;
// 	// logic [63:0] tb_input_test_370 = 64'h94d78cf57cd6e7ea;
// 	// logic [63:0] tb_input_test_371 = 64'ha6b6550f8249ec6b;
// 	// logic [63:0] tb_input_test_372 = 64'hc19ae84ef27de757;
// 	// logic [63:0] tb_input_test_373 = 64'he2557ade0747e253;
// 	// logic [63:0] tb_input_test_374 = 64'hc0282fdd809932d6;
// 	// logic [63:0] tb_input_test_375 = 64'hd3fbb2bdab97dc48;
// 	// logic [63:0] tb_input_test_376 = 64'had21d99d7daabf2f;
// 	// logic [63:0] tb_input_test_377 = 64'h982adc6f0d3c26b3;
// 	// logic [63:0] tb_input_test_378 = 64'h95e9a3d4d09dd034;
// 	// logic [63:0] tb_input_test_379 = 64'ha2a61b7e14e8816f;
// 	// logic [63:0] tb_input_test_380 = 64'hf422d9fb362f6b12;
// 	// logic [63:0] tb_input_test_381 = 64'h98c1c847508f2ccf;
// 	// logic [63:0] tb_input_test_382 = 64'heb1f31a257e38e72;
// 	// logic [63:0] tb_input_test_383 = 64'hfd7eabbe442991f1;
// 	// logic [63:0] tb_input_test_384 = 64'hc23ef4cf143540f8;
// 	// logic [63:0] tb_input_test_385 = 64'h8069ba4e7c8d6b6b;
// 	// logic [63:0] tb_input_test_386 = 64'h9a26f238fb490a4a;
// 	// logic [63:0] tb_input_test_387 = 64'he447e533bbcfec17;
// 	// logic [63:0] tb_input_test_388 = 64'hc78189f862a33b04;
// 	// logic [63:0] tb_input_test_389 = 64'h8cb23ba93741cb68;
// 	// logic [63:0] tb_input_test_390 = 64'hd70aaf3c61459e8f;
// 	// logic [63:0] tb_input_test_391 = 64'h9d07b7b963a545e5;
// 	// logic [63:0] tb_input_test_392 = 64'h807693cb48bb734e;
// 	// logic [63:0] tb_input_test_393 = 64'hba49d606c90f9487;
// 	// logic [63:0] tb_input_test_394 = 64'h8606246c4cdce5a5;
// 	// logic [63:0] tb_input_test_395 = 64'hb3655b9a5b147943;
// 	// logic [63:0] tb_input_test_396 = 64'hc43edef9a91ac0a0;
// 	// logic [63:0] tb_input_test_397 = 64'hc3efcd7d97c6ac8e;
// 	// logic [63:0] tb_input_test_398 = 64'hf3288e08b6fd3006;
// 	// logic [63:0] tb_input_test_399 = 64'hee5432266d23ba37;
// 	// logic [63:0] tb_input_test_400 = 64'hcdcfe247d456f0bf;
// 	// logic [63:0] tb_input_test_401 = 64'ha3aef4062845b864;
// 	// logic [63:0] tb_input_test_402 = 64'he9ecccc864a90482;
// 	// logic [63:0] tb_input_test_403 = 64'hceed93b63dd377af;
// 	// logic [63:0] tb_input_test_404 = 64'h91859fcb30f4ae20;
// 	// logic [63:0] tb_input_test_405 = 64'hc46bf4721d29c4ee;
// 	// logic [63:0] tb_input_test_406 = 64'he6892fe44fb09e0d;
// 	// logic [63:0] tb_input_test_407 = 64'hb787b926fb0870b6;
// 	// logic [63:0] tb_input_test_408 = 64'hcd220b1205d6558c;
// 	// logic [63:0] tb_input_test_409 = 64'hd96c378d44697ac7;
// 	// logic [63:0] tb_input_test_410 = 64'ha423ae9b4028dae1;
// 	// logic [63:0] tb_input_test_411 = 64'he2ff65bed1381c59;
// 	// logic [63:0] tb_input_test_412 = 64'h880f3af012789f10;
// 	// logic [63:0] tb_input_test_413 = 64'hd3b89cb0c38a2148;
// 	// logic [63:0] tb_input_test_414 = 64'h9c907a058d19c5c3;
// 	// logic [63:0] tb_input_test_415 = 64'hb9147b31bf3cdb69;
// 	// logic [63:0] tb_input_test_416 = 64'h836f0aefce0c3023;
// 	// logic [63:0] tb_input_test_417 = 64'h89409fcf2515fbed;
// 	// logic [63:0] tb_input_test_418 = 64'h94a57945c7a08570;
// 	// logic [63:0] tb_input_test_419 = 64'hb3e26d44c725ce14;
// 	// logic [63:0] tb_input_test_420 = 64'h9d0cd56bb2db0126;
// 	// logic [63:0] tb_input_test_421 = 64'hd11e97b65c2bff8a;
// 	// logic [63:0] tb_input_test_422 = 64'hb3bd305be424e575;
// 	// logic [63:0] tb_input_test_423 = 64'hd3f23f651e477634;
// 	// logic [63:0] tb_input_test_424 = 64'hdd1475b304ed5ea2;
// 	// logic [63:0] tb_input_test_425 = 64'hbd51cae0a2e7494a;
// 	// logic [63:0] tb_input_test_426 = 64'hdff7611a0b153725;
// 	// logic [63:0] tb_input_test_427 = 64'hbb4a3abbacc908fe;
// 	// logic [63:0] tb_input_test_428 = 64'hfe88a167e9c02be7;
// 	// logic [63:0] tb_input_test_429 = 64'he646ec704aa5aeb8;
// 	// logic [63:0] tb_input_test_430 = 64'h8f9b1ba14c220915;
// 	// logic [63:0] tb_input_test_431 = 64'hac681f6e5226f758;
// 	// logic [63:0] tb_input_test_432 = 64'he8d4a452a86329b2;
// 	// logic [63:0] tb_input_test_433 = 64'h82987b17f6281777;
// 	// logic [63:0] tb_input_test_434 = 64'hf3f8d5fd16deb533;
// 	// logic [63:0] tb_input_test_435 = 64'h96f25d6fa0e4d4ec;
// 	// logic [63:0] tb_input_test_436 = 64'h8db67bac915bc545;
// 	// logic [63:0] tb_input_test_437 = 64'hcb3c3c6028e4686e;
// 	// logic [63:0] tb_input_test_438 = 64'hcf7e9f1e49f5c611;
// 	// logic [63:0] tb_input_test_439 = 64'hd9fbf7324e50f33e;
// 	// logic [63:0] tb_input_test_440 = 64'hac3ade60313a5c8e;
// 	// logic [63:0] tb_input_test_441 = 64'hbc30b6da8012e5b2;
// 	// logic [63:0] tb_input_test_442 = 64'h9fd5f94ba18ed511;
// 	// logic [63:0] tb_input_test_443 = 64'hbde5a44d5ce71901;
// 	// logic [63:0] tb_input_test_444 = 64'h8b6f52b6f9f81c0f;
// 	// logic [63:0] tb_input_test_445 = 64'haad3cb45ab7fcfd0;
// 	// logic [63:0] tb_input_test_446 = 64'hc68a73c1a24b6671;
// 	// logic [63:0] tb_input_test_447 = 64'ha66609763b53b2df;
// 	// logic [63:0] tb_input_test_448 = 64'hef8ace7b9b4425b6;
// 	// logic [63:0] tb_input_test_449 = 64'h87c3426e10ebc02f;
// 	// logic [63:0] tb_input_test_450 = 64'he236d2a74ab66f46;
// 	// logic [63:0] tb_input_test_451 = 64'hc955b66007759547;
// 	// logic [63:0] tb_input_test_452 = 64'h99a67114aa7fb1b8;
// 	// logic [63:0] tb_input_test_453 = 64'hdd5c3f97954ff533;
// 	// logic [63:0] tb_input_test_454 = 64'ha6a330eec4542605;
// 	// logic [63:0] tb_input_test_455 = 64'ha821dc277d07bce9;
// 	// logic [63:0] tb_input_test_456 = 64'h9e544f47088a7aeb;
// 	// logic [63:0] tb_input_test_457 = 64'hb22719c7f8340c81;
// 	// logic [63:0] tb_input_test_458 = 64'h9d2b98d19cd64feb;
// 	// logic [63:0] tb_input_test_459 = 64'hefdb4cca542155b3;
// 	// logic [63:0] tb_input_test_460 = 64'heb467fe3a80ccee2;
// 	// logic [63:0] tb_input_test_461 = 64'h8309f6474fef631f;
// 	// logic [63:0] tb_input_test_462 = 64'h8afcf59802ea448e;
// 	// logic [63:0] tb_input_test_463 = 64'ha2002bb737a58901;
// 	// logic [63:0] tb_input_test_464 = 64'ha520c905d45dff8d;
// 	// logic [63:0] tb_input_test_465 = 64'hef5252879eca7aec;
// 	// logic [63:0] tb_input_test_466 = 64'hdc5429db575bc649;
// 	// logic [63:0] tb_input_test_467 = 64'hf5b2d103f73bd0d3;
// 	// logic [63:0] tb_input_test_468 = 64'h95135815485bed65;
// 	// logic [63:0] tb_input_test_469 = 64'hc1e43c6c2ea65ede;
// 	// logic [63:0] tb_input_test_470 = 64'hbe5e4cd2ad160246;
// 	// logic [63:0] tb_input_test_471 = 64'hdd45e8752a62493f;
// 	// logic [63:0] tb_input_test_472 = 64'he185615030d99a9c;
// 	// logic [63:0] tb_input_test_473 = 64'hcdb130e9487d878f;
// 	// logic [63:0] tb_input_test_474 = 64'hd1749d992b503c14;
// 	// logic [63:0] tb_input_test_475 = 64'hc1567a25fca5a0db;
// 	// logic [63:0] tb_input_test_476 = 64'hcca894da9d2c564b;
// 	// logic [63:0] tb_input_test_477 = 64'h96f42e5d246d4bbf;
// 	// logic [63:0] tb_input_test_478 = 64'hb9aa1ee15a6c6c79;
// 	// logic [63:0] tb_input_test_479 = 64'hfa14cbed74c73be1;
// 	// logic [63:0] tb_input_test_480 = 64'hf93158958300e5a9;
// 	// logic [63:0] tb_input_test_481 = 64'ha4b7055e95d2cb80;
// 	// logic [63:0] tb_input_test_482 = 64'hc5c31df3daa0a807;
// 	// logic [63:0] tb_input_test_483 = 64'haf8e9a32414f9d29;
// 	// logic [63:0] tb_input_test_484 = 64'hb35e8b13e65e45e1;
// 	// logic [63:0] tb_input_test_485 = 64'hdf19022e54467e88;
// 	// logic [63:0] tb_input_test_486 = 64'h9115f541eaea0e7a;
// 	// logic [63:0] tb_input_test_487 = 64'hf14b84ea7e9a1ca2;
// 	// logic [63:0] tb_input_test_488 = 64'hbc20998e44c629e1;
// 	// logic [63:0] tb_input_test_489 = 64'hd38af4bb57e5f1c1;
// 	// logic [63:0] tb_input_test_490 = 64'hb8ef48cadfa8cdc0;
// 	// logic [63:0] tb_input_test_491 = 64'hae051b671c7d1b5d;
// 	// logic [63:0] tb_input_test_492 = 64'he91afec691c99cb4;
// 	// logic [63:0] tb_input_test_493 = 64'he798ce3f46469365;
// 	// logic [63:0] tb_input_test_494 = 64'hafd3380fd8850f63;
// 	// logic [63:0] tb_input_test_495 = 64'h98dacc905ea52a04;
// 	// logic [63:0] tb_input_test_496 = 64'ha56ebf8e9d312460;
// 	// logic [63:0] tb_input_test_497 = 64'h9eda2938f387ffc8;
// 	// logic [63:0] tb_input_test_498 = 64'ha78904ea01263d6c;
// 	// logic [63:0] tb_input_test_499 = 64'h8d27d34d5cc23eba;


// // tb_input_block = tb_input_test_0;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_1;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_2;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_3;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_4;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_5;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_6;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_7;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_8;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_9;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_10;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_11;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_12;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_13;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_14;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_15;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_16;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_17;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_18;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_19;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_20;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_21;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_22;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_23;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_24;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_25;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_26;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_27;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_28;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_29;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_30;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_31;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_32;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_33;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_34;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_35;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_36;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_37;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_38;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_39;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_40;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_41;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_42;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_43;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_44;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_45;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_46;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_47;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_48;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_49;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_50;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_51;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_52;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_53;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_54;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_55;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_56;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_57;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_58;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_59;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_60;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_61;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_62;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_63;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_64;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_65;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_66;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_67;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_68;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_69;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_70;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_71;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_72;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_73;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_74;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_75;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_76;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_77;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_78;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_79;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_80;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_81;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_82;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_83;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_84;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_85;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_86;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_87;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_88;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_89;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_90;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_91;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_92;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_93;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_94;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_95;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_96;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_97;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_98;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_99;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_100;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_101;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_102;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_103;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_104;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_105;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_106;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_107;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_108;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_109;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_110;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_111;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_112;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_113;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_114;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_115;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_116;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_117;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_118;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_119;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_120;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_121;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_122;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_123;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_124;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_125;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_126;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_127;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_128;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_129;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_130;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_131;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_132;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_133;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_134;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_135;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_136;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_137;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_138;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_139;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_140;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_141;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_142;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_143;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_144;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_145;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_146;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_147;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_148;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_149;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_150;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_151;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_152;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_153;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_154;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_155;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_156;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_157;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_158;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_159;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_160;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_161;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_162;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_163;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_164;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_165;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_166;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_167;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_168;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_169;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_170;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_171;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_172;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_173;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_174;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_175;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_176;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_177;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_178;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_179;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_180;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_181;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_182;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_183;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_184;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_185;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_186;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_187;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_188;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_189;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_190;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_191;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_192;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_193;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_194;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_195;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_196;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_197;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_198;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_199;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_200;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_201;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_202;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_203;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_204;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_205;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_206;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_207;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_208;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_209;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_210;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_211;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_212;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_213;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_214;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_215;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_216;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_217;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_218;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_219;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_220;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_221;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_222;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_223;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_224;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_225;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_226;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_227;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_228;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_229;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_230;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_231;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_232;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_233;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_234;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_235;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_236;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_237;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_238;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_239;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_240;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_241;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_242;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_243;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_244;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_245;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_246;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_247;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_248;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_249;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_250;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_251;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_252;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_253;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_254;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_255;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_256;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_257;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_258;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_259;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_260;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_261;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_262;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_263;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_264;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_265;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_266;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_267;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_268;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_269;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_270;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_271;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_272;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_273;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_274;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_275;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_276;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_277;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_278;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_279;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_280;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_281;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_282;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_283;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_284;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_285;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_286;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_287;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_288;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_289;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_290;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_291;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_292;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_293;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_294;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_295;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_296;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_297;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_298;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_299;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_300;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_301;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_302;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_303;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_304;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_305;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_306;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_307;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_308;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_309;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_310;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_311;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_312;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_313;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_314;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_315;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_316;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_317;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_318;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_319;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_320;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_321;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_322;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_323;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_324;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_325;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_326;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_327;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_328;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_329;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_330;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_331;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_332;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_333;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_334;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_335;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_336;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_337;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_338;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_339;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_340;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_341;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_342;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_343;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_344;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_345;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_346;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_347;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_348;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_349;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_350;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_351;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_352;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_353;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_354;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_355;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_356;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_357;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_358;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_359;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_360;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_361;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_362;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_363;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_364;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_365;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_366;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_367;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_368;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_369;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_370;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_371;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_372;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_373;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_374;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_375;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_376;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_377;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_378;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_379;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_380;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_381;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_382;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_383;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_384;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_385;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_386;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_387;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_388;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_389;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_390;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_391;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_392;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_393;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_394;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_395;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_396;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_397;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_398;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_399;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_400;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_401;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_402;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_403;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_404;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_405;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_406;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_407;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_408;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_409;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_410;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_411;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_412;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_413;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_414;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_415;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_416;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_417;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_418;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_419;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_420;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_421;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_422;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_423;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_424;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_425;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_426;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_427;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_428;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_429;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_430;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_431;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_432;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_433;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_434;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_435;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_436;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_437;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_438;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_439;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_440;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_441;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_442;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_443;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_444;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_445;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_446;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_447;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_448;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_449;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_450;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_451;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_452;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_453;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_454;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_455;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_456;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_457;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_458;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_459;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_460;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_461;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_462;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_463;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_464;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_465;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_466;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_467;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_468;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_469;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_470;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_471;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_472;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_473;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_474;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_475;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_476;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_477;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_478;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_479;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_480;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_481;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_482;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_483;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_484;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_485;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_486;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_487;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_488;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_489;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_490;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_491;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_492;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_493;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_494;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_495;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_496;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_497;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_498;

// // @(negedge tb_clk);
// // tb_input_block = tb_input_test_499;


// //	end


// endmodule
